library verilog;
use verilog.vl_types.all;
entity tagArray is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        we              : in     vl_logic_vector(127 downto 0);
        tag             : in     vl_logic_vector(6 downto 0);
        tagOut0         : out    vl_logic_vector(5 downto 0);
        tagOut1         : out    vl_logic_vector(5 downto 0);
        tagOut2         : out    vl_logic_vector(5 downto 0);
        tagOut3         : out    vl_logic_vector(5 downto 0);
        tagOut4         : out    vl_logic_vector(5 downto 0);
        tagOut5         : out    vl_logic_vector(5 downto 0);
        tagOut6         : out    vl_logic_vector(5 downto 0);
        tagOut7         : out    vl_logic_vector(5 downto 0);
        tagOut8         : out    vl_logic_vector(5 downto 0);
        tagOut9         : out    vl_logic_vector(5 downto 0);
        tagOut10        : out    vl_logic_vector(5 downto 0);
        tagOut11        : out    vl_logic_vector(5 downto 0);
        tagOut12        : out    vl_logic_vector(5 downto 0);
        tagOut13        : out    vl_logic_vector(5 downto 0);
        tagOut14        : out    vl_logic_vector(5 downto 0);
        tagOut15        : out    vl_logic_vector(5 downto 0);
        tagOut16        : out    vl_logic_vector(5 downto 0);
        tagOut17        : out    vl_logic_vector(5 downto 0);
        tagOut18        : out    vl_logic_vector(5 downto 0);
        tagOut19        : out    vl_logic_vector(5 downto 0);
        tagOut20        : out    vl_logic_vector(5 downto 0);
        tagOut21        : out    vl_logic_vector(5 downto 0);
        tagOut22        : out    vl_logic_vector(5 downto 0);
        tagOut23        : out    vl_logic_vector(5 downto 0);
        tagOut24        : out    vl_logic_vector(5 downto 0);
        tagOut25        : out    vl_logic_vector(5 downto 0);
        tagOut26        : out    vl_logic_vector(5 downto 0);
        tagOut27        : out    vl_logic_vector(5 downto 0);
        tagOut28        : out    vl_logic_vector(5 downto 0);
        tagOut29        : out    vl_logic_vector(5 downto 0);
        tagOut30        : out    vl_logic_vector(5 downto 0);
        tagOut31        : out    vl_logic_vector(5 downto 0);
        tagOut32        : out    vl_logic_vector(5 downto 0);
        tagOut33        : out    vl_logic_vector(5 downto 0);
        tagOut34        : out    vl_logic_vector(5 downto 0);
        tagOut35        : out    vl_logic_vector(5 downto 0);
        tagOut36        : out    vl_logic_vector(5 downto 0);
        tagOut37        : out    vl_logic_vector(5 downto 0);
        tagOut38        : out    vl_logic_vector(5 downto 0);
        tagOut39        : out    vl_logic_vector(5 downto 0);
        tagOut40        : out    vl_logic_vector(5 downto 0);
        tagOut41        : out    vl_logic_vector(5 downto 0);
        tagOut42        : out    vl_logic_vector(5 downto 0);
        tagOut43        : out    vl_logic_vector(5 downto 0);
        tagOut44        : out    vl_logic_vector(5 downto 0);
        tagOut45        : out    vl_logic_vector(5 downto 0);
        tagOut46        : out    vl_logic_vector(5 downto 0);
        tagOut47        : out    vl_logic_vector(5 downto 0);
        tagOut48        : out    vl_logic_vector(5 downto 0);
        tagOut49        : out    vl_logic_vector(5 downto 0);
        tagOut50        : out    vl_logic_vector(5 downto 0);
        tagOut51        : out    vl_logic_vector(5 downto 0);
        tagOut52        : out    vl_logic_vector(5 downto 0);
        tagOut53        : out    vl_logic_vector(5 downto 0);
        tagOut54        : out    vl_logic_vector(5 downto 0);
        tagOut55        : out    vl_logic_vector(5 downto 0);
        tagOut56        : out    vl_logic_vector(5 downto 0);
        tagOut57        : out    vl_logic_vector(5 downto 0);
        tagOut58        : out    vl_logic_vector(5 downto 0);
        tagOut59        : out    vl_logic_vector(5 downto 0);
        tagOut60        : out    vl_logic_vector(5 downto 0);
        tagOut61        : out    vl_logic_vector(5 downto 0);
        tagOut62        : out    vl_logic_vector(5 downto 0);
        tagOut63        : out    vl_logic_vector(5 downto 0);
        tagOut64        : out    vl_logic_vector(5 downto 0);
        tagOut65        : out    vl_logic_vector(5 downto 0);
        tagOut66        : out    vl_logic_vector(5 downto 0);
        tagOut67        : out    vl_logic_vector(5 downto 0);
        tagOut68        : out    vl_logic_vector(5 downto 0);
        tagOut69        : out    vl_logic_vector(5 downto 0);
        tagOut70        : out    vl_logic_vector(5 downto 0);
        tagOut71        : out    vl_logic_vector(5 downto 0);
        tagOut72        : out    vl_logic_vector(5 downto 0);
        tagOut73        : out    vl_logic_vector(5 downto 0);
        tagOut74        : out    vl_logic_vector(5 downto 0);
        tagOut75        : out    vl_logic_vector(5 downto 0);
        tagOut76        : out    vl_logic_vector(5 downto 0);
        tagOut77        : out    vl_logic_vector(5 downto 0);
        tagOut78        : out    vl_logic_vector(5 downto 0);
        tagOut79        : out    vl_logic_vector(5 downto 0);
        tagOut80        : out    vl_logic_vector(5 downto 0);
        tagOut81        : out    vl_logic_vector(5 downto 0);
        tagOut82        : out    vl_logic_vector(5 downto 0);
        tagOut83        : out    vl_logic_vector(5 downto 0);
        tagOut84        : out    vl_logic_vector(5 downto 0);
        tagOut85        : out    vl_logic_vector(5 downto 0);
        tagOut86        : out    vl_logic_vector(5 downto 0);
        tagOut87        : out    vl_logic_vector(5 downto 0);
        tagOut88        : out    vl_logic_vector(5 downto 0);
        tagOut89        : out    vl_logic_vector(5 downto 0);
        tagOut90        : out    vl_logic_vector(5 downto 0);
        tagOut91        : out    vl_logic_vector(5 downto 0);
        tagOut92        : out    vl_logic_vector(5 downto 0);
        tagOut93        : out    vl_logic_vector(5 downto 0);
        tagOut94        : out    vl_logic_vector(5 downto 0);
        tagOut95        : out    vl_logic_vector(5 downto 0);
        tagOut96        : out    vl_logic_vector(5 downto 0);
        tagOut97        : out    vl_logic_vector(5 downto 0);
        tagOut98        : out    vl_logic_vector(5 downto 0);
        tagOut99        : out    vl_logic_vector(5 downto 0);
        tagOut100       : out    vl_logic_vector(5 downto 0);
        tagOut101       : out    vl_logic_vector(5 downto 0);
        tagOut102       : out    vl_logic_vector(5 downto 0);
        tagOut103       : out    vl_logic_vector(5 downto 0);
        tagOut104       : out    vl_logic_vector(5 downto 0);
        tagOut105       : out    vl_logic_vector(5 downto 0);
        tagOut106       : out    vl_logic_vector(5 downto 0);
        tagOut107       : out    vl_logic_vector(5 downto 0);
        tagOut108       : out    vl_logic_vector(5 downto 0);
        tagOut109       : out    vl_logic_vector(5 downto 0);
        tagOut110       : out    vl_logic_vector(5 downto 0);
        tagOut111       : out    vl_logic_vector(5 downto 0);
        tagOut112       : out    vl_logic_vector(5 downto 0);
        tagOut113       : out    vl_logic_vector(5 downto 0);
        tagOut114       : out    vl_logic_vector(5 downto 0);
        tagOut115       : out    vl_logic_vector(5 downto 0);
        tagOut116       : out    vl_logic_vector(5 downto 0);
        tagOut117       : out    vl_logic_vector(5 downto 0);
        tagOut118       : out    vl_logic_vector(5 downto 0);
        tagOut119       : out    vl_logic_vector(5 downto 0);
        tagOut120       : out    vl_logic_vector(5 downto 0);
        tagOut121       : out    vl_logic_vector(5 downto 0);
        tagOut122       : out    vl_logic_vector(5 downto 0);
        tagOut123       : out    vl_logic_vector(5 downto 0);
        tagOut124       : out    vl_logic_vector(5 downto 0);
        tagOut125       : out    vl_logic_vector(5 downto 0);
        tagOut126       : out    vl_logic_vector(5 downto 0);
        tagOut127       : out    vl_logic_vector(5 downto 0)
    );
end tagArray;
