library verilog;
use verilog.vl_types.all;
entity processorKiTestBench is
end processorKiTestBench;
